---------------------------------------------------------------------------
-- Company     : Universidade Federal de Santa Catarina
-- Author(s)   : Victor H B Preuss
--
-- Creation Date : 12/04/2018
-- File          : rom.vhd
--
-- Abstract :
--
---------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;

---------------------------------------------------------------------------
entity rom is
    generic (
        DATA_SIZE   : integer := 16; -- size of an addressable data
        ADDR_SIZE   : integer := 10; -- number of bits of and address
        MEM_SIZE    : integer := 1024 -- memory size
    );
    port (
        addr    : in std_logic_vector(ADDR_SIZE-1 downto 0);
        data    : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
end entity;

---------------------------------------------------------------------------
architecture arch of rom is

    subtype word_t is std_logic_vector(DATA_SIZE-1 downto 0);
    type memory_t is array(0 to MEM_SIZE-1) of word_t;

    --signal addr_reg : integer := 0;
    signal addri : integer := 0;
    constant rom_data : memory_t := (
				x"310D",
				x"320E",
				x"F410",
				x"F420",
				x"F410",
				x"F420",
				x"F510",
				x"F520",
				x"F410",
				x"F420",
				x"F800",
				x"F801",
				x"F800",
				x"F801",
				x"F800",
				x"F801",
				x"F901",
				x"F900",
				x"F050",
				x"F050",
				x"F050",
				x"F050",
				x"F050",
				x"F060",
				x"F060",
				x"F060",
				x"F060",
				x"F060",
				x"F150",
				x"F150",
				x"F160",
				x"F901",
				x"F900",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF");

begin

    addri <= to_integer(unsigned(addr));
    data <= rom_data(addri);

end architecture;