---------------------------------------------------------------------------
-- Company     : Universidade Federal de Santa Catarina
-- Author(s)   : Victor H B Preuss
--
-- Creation Date : 12/04/2018
-- File          : rom.vhd
--
-- Abstract :
--
---------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;

---------------------------------------------------------------------------
entity rom is
    generic (
        DATA_SIZE   : integer := 16; -- size of an addressable data
        ADDR_SIZE   : integer := 10; -- number of bits of and address
        MEM_SIZE    : integer := 1024 -- memory size
    );
    port (
        addr    : in std_logic_vector(ADDR_SIZE-1 downto 0);
        data    : out std_logic_vector(DATA_SIZE-1 downto 0)
    );
end entity;

---------------------------------------------------------------------------
architecture arch of rom is

    subtype word_t is std_logic_vector(DATA_SIZE-1 downto 0);
    type memory_t is array(0 to MEM_SIZE-1) of word_t;

    --signal addr_reg : integer := 0;
    signal addri : integer := 0;
    constant rom_data : memory_t := (
				x"D309",
				x"D804",
				x"D303",
				x"D805",
				x"D306",
				x"D806",
				x"D302",
				x"D807",
				x"D308",
				x"D808",
				x"D301",
				x"D809",
				x"D304",
				x"D80A",
				x"D305",
				x"D80B",
				x"2823",
				x"D313",
				x"D804",
				x"D30D",
				x"D805",
				x"D310",
				x"D806",
				x"D30C",
				x"D807",
				x"D312",
				x"D808",
				x"D30B",
				x"D809",
				x"D30E",
				x"D80A",
				x"D30F",
				x"D80B",
				x"2823",
				x"0800",
				x"D000",
				x"D301",
				x"D802",
				x"3200",
				x"D202",
				x"D030",
				x"D308",
				x"7003",
				x"182F",
				x"142E",
				x"102F",
				x"3201",
				x"E46F",
				x"D300",
				x"D803",
				x"3300",
				x"D203",
				x"D040",
				x"D307",
				x"7004",
				x"183B",
				x"143A",
				x"103B",
				x"3301",
				x"E86D",
				x"3400",
				x"D203",
				x"D060",
				x"D006",
				x"8304",
				x"D150",
				x"D203",
				x"D070",
				x"D301",
				x"8070",
				x"D007",
				x"8304",
				x"D160",
				x"7056",
				x"184E",
				x"144D",
				x"104E",
				x"3401",
				x"EC6B",
				x"D203",
				x"D060",
				x"D006",
				x"8304",
				x"D150",
				x"D005",
				x"D80C",
				x"D203",
				x"D060",
				x"D301",
				x"8060",
				x"D006",
				x"8304",
				x"D150",
				x"D203",
				x"D060",
				x"D006",
				x"8304",
				x"D405",
				x"D20C",
				x"D050",
				x"D203",
				x"D060",
				x"D301",
				x"8060",
				x"D006",
				x"8304",
				x"D405",
				x"F803",
				x"0832",
				x"F802",
				x"0826",
				x"3080",
				x"D380",
				x"DC1A",
				x"0872",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF",
				x"FFFF");

begin

    addri <= to_integer(unsigned(addr));
    data <= rom_data(addri);

end architecture;